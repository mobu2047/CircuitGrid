.title Active DC Circuit
R 0 1 73m
R 3 1 65
R 0 2 98m
I 2 3 18


.control
op
.endc
.end
