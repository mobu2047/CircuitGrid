.title Active DC Circuit
R 0 1 73m
R 3 1 65
R 0 2 5m
I 2 3 94


.control
op
.endc
.end
