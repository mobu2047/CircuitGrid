.title Active DC Circuit
.MODEL NPN_MODEL NPN
R 19 20 0
V 19 28 0
R 12 29 0
V 29 28 0
QT 28 20 12 NPN_MODEL


.control
op
.endc
.end
