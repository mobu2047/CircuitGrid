.title Active DC Circuit
R 24 25 0
V 24 32 0


.control
op
.endc
.end
