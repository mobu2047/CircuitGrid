.title Active DC Circuit
R3 1 0 <Empty>
I1 2 0 <Empty>
R1 3 1 <Empty>
R2 4 2 <Empty>
R4 4 3 <Empty>


.control
op
print v(2, 4) ; measurement of U1
.endc
.end
