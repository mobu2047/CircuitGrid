.title Active DC Circuit
E2 0 1 0 2 <Empty>
R1 0 2 <Empty>
E1 1 2 0 2 <Empty>
I1 3 2 <Empty>
I2 2 4 <Empty>
I3 4 3 <Empty>
R2 4 3 <Empty>


.control
op
print -v(2) ; measurement of U0
.endc
.end
