.title Active DC Circuit
R 0 1 58
R 2 1 65
R 4 1 84
R 3 2 51
R 0 4 66
I 2 4 60
R 3 2 24


.control
op
print -v(1) ; measurement of U0
.endc
.end
