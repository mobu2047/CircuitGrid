.title Active DC Circuit
R 0 1 29k
R 2 0 500k
R 3 1 2k
R 2 3 52
R 2 4 28
V 4 3 33


.control
op
.endc
.end
